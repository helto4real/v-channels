
module channel

pub struct Channel {

}